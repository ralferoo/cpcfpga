-- bootrom.vhd
library IEEE;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.std_logic_arith.all;

entity bootrom is
    port(
	clk		: in  std_logic;
        addr		: in  std_logic_vector(13 downto 0);
        data		: out std_logic_vector(7 downto 0)
    );
end bootrom;

architecture impl of bootrom is


begin


process (addr)
    begin

	        case addr(9 downto 0) is 
                    when "0000000000" => data <= X"f3";
                    when "0000000001" => data <= X"31";
                    when "0000000010" => data <= X"fe";
                    when "0000000011" => data <= X"bf";
                    when "0000000100" => data <= X"01";
                    when "0000000101" => data <= X"8d";
                    when "0000000110" => data <= X"7f";
                    when "0000000111" => data <= X"ed";
                    when "0000001000" => data <= X"49";
                    when "0000001001" => data <= X"01";
                    when "0000001010" => data <= X"de";
                    when "0000001011" => data <= X"fa";
                    when "0000001100" => data <= X"ed";
                    when "0000001101" => data <= X"78";
                    when "0000001110" => data <= X"0b";
                    when "0000001111" => data <= X"e6";
                    when "0000010000" => data <= X"01";
                    when "0000010001" => data <= X"ca";
                    when "0000010010" => data <= X"b2";
                    when "0000010011" => data <= X"01";
                    when "0000010100" => data <= X"01";
                    when "0000010101" => data <= X"dd";
                    when "0000010110" => data <= X"fa";
                    when "0000010111" => data <= X"dd";
                    when "0000011000" => data <= X"26";
                    when "0000011001" => data <= X"80";
                    when "0000011010" => data <= X"21";
                    when "0000011011" => data <= X"68";
                    when "0000011100" => data <= X"01";
                    when "0000011101" => data <= X"cd";
                    when "0000011110" => data <= X"f4";
                    when "0000011111" => data <= X"00";
                    when "0000100000" => data <= X"cd";
                    when "0000100001" => data <= X"2a";
                    when "0000100010" => data <= X"01";
                    when "0000100011" => data <= X"fe";
                    when "0000100100" => data <= X"53";
                    when "0000100101" => data <= X"28";
                    when "0000100110" => data <= X"14";
                    when "0000100111" => data <= X"fe";
                    when "0000101000" => data <= X"0d";
                    when "0000101001" => data <= X"28";
                    when "0000101010" => data <= X"09";
                    when "0000101011" => data <= X"fe";
                    when "0000101100" => data <= X"0a";
                    when "0000101101" => data <= X"28";
                    when "0000101110" => data <= X"05";
                    when "0000101111" => data <= X"cd";
                    when "0000110000" => data <= X"2a";
                    when "0000110001" => data <= X"01";
                    when "0000110010" => data <= X"18";
                    when "0000110011" => data <= X"ef";
                    when "0000110100" => data <= X"cd";
                    when "0000110101" => data <= X"2a";
                    when "0000110110" => data <= X"01";
                    when "0000110111" => data <= X"fe";
                    when "0000111000" => data <= X"53";
                    when "0000111001" => data <= X"20";
                    when "0000111010" => data <= X"e8";
                    when "0000111011" => data <= X"cd";
                    when "0000111100" => data <= X"2a";
                    when "0000111101" => data <= X"01";
                    when "0000111110" => data <= X"fe";
                    when "0000111111" => data <= X"30";
                    when "0001000000" => data <= X"28";
                    when "0001000001" => data <= X"2a";
                    when "0001000010" => data <= X"fe";
                    when "0001000011" => data <= X"31";
                    when "0001000100" => data <= X"28";
                    when "0001000101" => data <= X"48";
                    when "0001000110" => data <= X"fe";
                    when "0001000111" => data <= X"35";
                    when "0001001000" => data <= X"28";
                    when "0001001001" => data <= X"64";
                    when "0001001010" => data <= X"fe";
                    when "0001001011" => data <= X"39";
                    when "0001001100" => data <= X"20";
                    when "0001001101" => data <= X"7f";
                    when "0001001110" => data <= X"cd";
                    when "0001001111" => data <= X"df";
                    when "0001010000" => data <= X"00";
                    when "0001010001" => data <= X"cd";
                    when "0001010010" => data <= X"be";
                    when "0001010011" => data <= X"00";
                    when "0001010100" => data <= X"e5";
                    when "0001010101" => data <= X"21";
                    when "0001010110" => data <= X"9a";
                    when "0001010111" => data <= X"01";
                    when "0001011000" => data <= X"cd";
                    when "0001011001" => data <= X"f4";
                    when "0001011010" => data <= X"00";
                    when "0001011011" => data <= X"e1";
                    when "0001011100" => data <= X"e5";
                    when "0001011101" => data <= X"7c";
                    when "0001011110" => data <= X"cd";
                    when "0001011111" => data <= X"03";
                    when "0001100000" => data <= X"01";
                    when "0001100001" => data <= X"7d";
                    when "0001100010" => data <= X"cd";
                    when "0001100011" => data <= X"03";
                    when "0001100100" => data <= X"01";
                    when "0001100101" => data <= X"21";
                    when "0001100110" => data <= X"97";
                    when "0001100111" => data <= X"01";
                    when "0001101000" => data <= X"cd";
                    when "0001101001" => data <= X"f4";
                    when "0001101010" => data <= X"00";
                    when "0001101011" => data <= X"c9";
                    when "0001101100" => data <= X"dd";
                    when "0001101101" => data <= X"21";
                    when "0001101110" => data <= X"00";
                    when "0001101111" => data <= X"00";
                    when "0001110000" => data <= X"cd";
                    when "0001110001" => data <= X"df";
                    when "0001110010" => data <= X"00";
                    when "0001110011" => data <= X"af";
                    when "0001110100" => data <= X"fd";
                    when "0001110101" => data <= X"b4";
                    when "0001110110" => data <= X"28";
                    when "0001110111" => data <= X"0b";
                    when "0001111000" => data <= X"cd";
                    when "0001111001" => data <= X"35";
                    when "0001111010" => data <= X"01";
                    when "0001111011" => data <= X"fd";
                    when "0001111100" => data <= X"25";
                    when "0001111101" => data <= X"0d";
                    when "0001111110" => data <= X"ed";
                    when "0001111111" => data <= X"79";
                    when "0010000000" => data <= X"0c";
                    when "0010000001" => data <= X"18";
                    when "0010000010" => data <= X"f0";
                    when "0010000011" => data <= X"cd";
                    when "0010000100" => data <= X"be";
                    when "0010000101" => data <= X"00";
                    when "0010000110" => data <= X"3e";
                    when "0010000111" => data <= X"20";
                    when "0010001000" => data <= X"0d";
                    when "0010001001" => data <= X"ed";
                    when "0010001010" => data <= X"79";
                    when "0010001011" => data <= X"0c";
                    when "0010001100" => data <= X"18";
                    when "0010001101" => data <= X"92";
                    when "0010001110" => data <= X"dd";
                    when "0010001111" => data <= X"7c";
                    when "0010010000" => data <= X"e6";
                    when "0010010001" => data <= X"80";
                    when "0010010010" => data <= X"20";
                    when "0010010011" => data <= X"8f";
                    when "0010010100" => data <= X"cd";
                    when "0010010101" => data <= X"df";
                    when "0010010110" => data <= X"00";
                    when "0010010111" => data <= X"af";
                    when "0010011000" => data <= X"fd";
                    when "0010011001" => data <= X"b4";
                    when "0010011010" => data <= X"28";
                    when "0010011011" => data <= X"09";
                    when "0010011100" => data <= X"cd";
                    when "0010011101" => data <= X"35";
                    when "0010011110" => data <= X"01";
                    when "0010011111" => data <= X"fd";
                    when "0010100000" => data <= X"25";
                    when "0010100001" => data <= X"77";
                    when "0010100010" => data <= X"23";
                    when "0010100011" => data <= X"18";
                    when "0010100100" => data <= X"f2";
                    when "0010100101" => data <= X"cd";
                    when "0010100110" => data <= X"be";
                    when "0010100111" => data <= X"00";
                    when "0010101000" => data <= X"dd";
                    when "0010101001" => data <= X"23";
                    when "0010101010" => data <= X"3e";
                    when "0010101011" => data <= X"2e";
                    when "0010101100" => data <= X"18";
                    when "0010101101" => data <= X"da";
                    when "0010101110" => data <= X"cd";
                    when "0010101111" => data <= X"df";
                    when "0010110000" => data <= X"00";
                    when "0010110001" => data <= X"cd";
                    when "0010110010" => data <= X"be";
                    when "0010110011" => data <= X"00";
                    when "0010110100" => data <= X"dd";
                    when "0010110101" => data <= X"e5";
                    when "0010110110" => data <= X"d1";
                    when "0010110111" => data <= X"a7";
                    when "0010111000" => data <= X"ed";
                    when "0010111001" => data <= X"52";
                    when "0010111010" => data <= X"28";
                    when "0010111011" => data <= X"d0";
                    when "0010111100" => data <= X"18";
                    when "0010111101" => data <= X"0f";
                    when "0010111110" => data <= X"cd";
                    when "0010111111" => data <= X"35";
                    when "0011000000" => data <= X"01";
                    when "0011000001" => data <= X"dd";
                    when "0011000010" => data <= X"7c";
                    when "0011000011" => data <= X"e6";
                    when "0011000100" => data <= X"80";
                    when "0011000101" => data <= X"20";
                    when "0011000110" => data <= X"c5";
                    when "0011000111" => data <= X"fd";
                    when "0011001000" => data <= X"7d";
                    when "0011001001" => data <= X"3c";
                    when "0011001010" => data <= X"fd";
                    when "0011001011" => data <= X"b4";
                    when "0011001100" => data <= X"c8";
                    when "0011001101" => data <= X"e1";
                    when "0011001110" => data <= X"dd";
                    when "0011001111" => data <= X"7c";
                    when "0011010000" => data <= X"e6";
                    when "0011010001" => data <= X"80";
                    when "0011010010" => data <= X"20";
                    when "0011010011" => data <= X"b8";
                    when "0011010100" => data <= X"dd";
                    when "0011010101" => data <= X"26";
                    when "0011010110" => data <= X"80";
                    when "0011010111" => data <= X"21";
                    when "0011011000" => data <= X"a8";
                    when "0011011001" => data <= X"01";
                    when "0011011010" => data <= X"cd";
                    when "0011011011" => data <= X"f4";
                    when "0011011100" => data <= X"00";
                    when "0011011101" => data <= X"18";
                    when "0011011110" => data <= X"ad";
                    when "0011011111" => data <= X"fd";
                    when "0011100000" => data <= X"2e";
                    when "0011100001" => data <= X"00";
                    when "0011100010" => data <= X"cd";
                    when "0011100011" => data <= X"35";
                    when "0011100100" => data <= X"01";
                    when "0011100101" => data <= X"d6";
                    when "0011100110" => data <= X"03";
                    when "0011100111" => data <= X"fd";
                    when "0011101000" => data <= X"67";
                    when "0011101001" => data <= X"38";
                    when "0011101010" => data <= X"e2";
                    when "0011101011" => data <= X"cd";
                    when "0011101100" => data <= X"35";
                    when "0011101101" => data <= X"01";
                    when "0011101110" => data <= X"67";
                    when "0011101111" => data <= X"cd";
                    when "0011110000" => data <= X"35";
                    when "0011110001" => data <= X"01";
                    when "0011110010" => data <= X"6f";
                    when "0011110011" => data <= X"c9";
                    when "0011110100" => data <= X"ed";
                    when "0011110101" => data <= X"78";
                    when "0011110110" => data <= X"17";
                    when "0011110111" => data <= X"30";
                    when "0011111000" => data <= X"fb";
                    when "0011111001" => data <= X"7e";
                    when "0011111010" => data <= X"b7";
                    when "0011111011" => data <= X"c8";
                    when "0011111100" => data <= X"0d";
                    when "0011111101" => data <= X"ed";
                    when "0011111110" => data <= X"79";
                    when "0011111111" => data <= X"0c";
                    when "0100000000" => data <= X"23";
                    when "0100000001" => data <= X"18";
                    when "0100000010" => data <= X"f1";
                    when "0100000011" => data <= X"f5";
                    when "0100000100" => data <= X"1f";
                    when "0100000101" => data <= X"1f";
                    when "0100000110" => data <= X"1f";
                    when "0100000111" => data <= X"1f";
                    when "0100001000" => data <= X"e6";
                    when "0100001001" => data <= X"0f";
                    when "0100001010" => data <= X"fe";
                    when "0100001011" => data <= X"0a";
                    when "0100001100" => data <= X"de";
                    when "0100001101" => data <= X"69";
                    when "0100001110" => data <= X"27";
                    when "0100001111" => data <= X"ed";
                    when "0100010000" => data <= X"70";
                    when "0100010001" => data <= X"f2";
                    when "0100010010" => data <= X"0f";
                    when "0100010011" => data <= X"01";
                    when "0100010100" => data <= X"0d";
                    when "0100010101" => data <= X"ed";
                    when "0100010110" => data <= X"79";
                    when "0100010111" => data <= X"0c";
                    when "0100011000" => data <= X"f1";
                    when "0100011001" => data <= X"e6";
                    when "0100011010" => data <= X"0f";
                    when "0100011011" => data <= X"fe";
                    when "0100011100" => data <= X"0a";
                    when "0100011101" => data <= X"de";
                    when "0100011110" => data <= X"69";
                    when "0100011111" => data <= X"27";
                    when "0100100000" => data <= X"ed";
                    when "0100100001" => data <= X"70";
                    when "0100100010" => data <= X"f2";
                    when "0100100011" => data <= X"20";
                    when "0100100100" => data <= X"01";
                    when "0100100101" => data <= X"0d";
                    when "0100100110" => data <= X"ed";
                    when "0100100111" => data <= X"79";
                    when "0100101000" => data <= X"0c";
                    when "0100101001" => data <= X"c9";
                    when "0100101010" => data <= X"ed";
                    when "0100101011" => data <= X"78";
                    when "0100101100" => data <= X"e6";
                    when "0100101101" => data <= X"40";
                    when "0100101110" => data <= X"28";
                    when "0100101111" => data <= X"fa";
                    when "0100110000" => data <= X"0d";
                    when "0100110001" => data <= X"ed";
                    when "0100110010" => data <= X"78";
                    when "0100110011" => data <= X"0c";
                    when "0100110100" => data <= X"c9";
                    when "0100110101" => data <= X"ed";
                    when "0100110110" => data <= X"78";
                    when "0100110111" => data <= X"e6";
                    when "0100111000" => data <= X"40";
                    when "0100111001" => data <= X"28";
                    when "0100111010" => data <= X"fa";
                    when "0100111011" => data <= X"0d";
                    when "0100111100" => data <= X"ed";
                    when "0100111101" => data <= X"78";
                    when "0100111110" => data <= X"0c";
                    when "0100111111" => data <= X"57";
                    when "0101000000" => data <= X"c6";
                    when "0101000001" => data <= X"c0";
                    when "0101000010" => data <= X"9f";
                    when "0101000011" => data <= X"e6";
                    when "0101000100" => data <= X"09";
                    when "0101000101" => data <= X"82";
                    when "0101000110" => data <= X"e6";
                    when "0101000111" => data <= X"0f";
                    when "0101001000" => data <= X"17";
                    when "0101001001" => data <= X"17";
                    when "0101001010" => data <= X"17";
                    when "0101001011" => data <= X"17";
                    when "0101001100" => data <= X"5f";
                    when "0101001101" => data <= X"ed";
                    when "0101001110" => data <= X"78";
                    when "0101001111" => data <= X"e6";
                    when "0101010000" => data <= X"40";
                    when "0101010001" => data <= X"28";
                    when "0101010010" => data <= X"fa";
                    when "0101010011" => data <= X"0d";
                    when "0101010100" => data <= X"ed";
                    when "0101010101" => data <= X"78";
                    when "0101010110" => data <= X"0c";
                    when "0101010111" => data <= X"57";
                    when "0101011000" => data <= X"c6";
                    when "0101011001" => data <= X"c0";
                    when "0101011010" => data <= X"9f";
                    when "0101011011" => data <= X"e6";
                    when "0101011100" => data <= X"09";
                    when "0101011101" => data <= X"82";
                    when "0101011110" => data <= X"e6";
                    when "0101011111" => data <= X"0f";
                    when "0101100000" => data <= X"b3";
                    when "0101100001" => data <= X"5f";
                    when "0101100010" => data <= X"fd";
                    when "0101100011" => data <= X"85";
                    when "0101100100" => data <= X"fd";
                    when "0101100101" => data <= X"6f";
                    when "0101100110" => data <= X"7b";
                    when "0101100111" => data <= X"c9";
                    when "0101101000" => data <= X"0d";
                    when "0101101001" => data <= X"0a";
                    when "0101101010" => data <= X"53";
                    when "0101101011" => data <= X"52";
                    when "0101101100" => data <= X"45";
                    when "0101101101" => data <= X"43";
                    when "0101101110" => data <= X"20";
                    when "0101101111" => data <= X"6c";
                    when "0101110000" => data <= X"6f";
                    when "0101110001" => data <= X"61";
                    when "0101110010" => data <= X"64";
                    when "0101110011" => data <= X"65";
                    when "0101110100" => data <= X"72";
                    when "0101110101" => data <= X"20";
                    when "0101110110" => data <= X"76";
                    when "0101110111" => data <= X"30";
                    when "0101111000" => data <= X"2e";
                    when "0101111001" => data <= X"30";
                    when "0101111010" => data <= X"32";
                    when "0101111011" => data <= X"62";
                    when "0101111100" => data <= X"2c";
                    when "0101111101" => data <= X"20";
                    when "0101111110" => data <= X"28";
                    when "0101111111" => data <= X"63";
                    when "0110000000" => data <= X"29";
                    when "0110000001" => data <= X"20";
                    when "0110000010" => data <= X"32";
                    when "0110000011" => data <= X"30";
                    when "0110000100" => data <= X"31";
                    when "0110000101" => data <= X"32";
                    when "0110000110" => data <= X"20";
                    when "0110000111" => data <= X"52";
                    when "0110001000" => data <= X"61";
                    when "0110001001" => data <= X"6e";
                    when "0110001010" => data <= X"75";
                    when "0110001011" => data <= X"6c";
                    when "0110001100" => data <= X"66";
                    when "0110001101" => data <= X"20";
                    when "0110001110" => data <= X"44";
                    when "0110001111" => data <= X"6f";
                    when "0110010000" => data <= X"73";
                    when "0110010001" => data <= X"77";
                    when "0110010010" => data <= X"65";
                    when "0110010011" => data <= X"6c";
                    when "0110010100" => data <= X"6c";
                    when "0110010101" => data <= X"0d";
                    when "0110010110" => data <= X"0a";
                    when "0110010111" => data <= X"0d";
                    when "0110011000" => data <= X"0a";
                    when "0110011001" => data <= X"00";
                    when "0110011010" => data <= X"0d";
                    when "0110011011" => data <= X"0a";
                    when "0110011100" => data <= X"4a";
                    when "0110011101" => data <= X"75";
                    when "0110011110" => data <= X"6d";
                    when "0110011111" => data <= X"70";
                    when "0110100000" => data <= X"69";
                    when "0110100001" => data <= X"6e";
                    when "0110100010" => data <= X"67";
                    when "0110100011" => data <= X"20";
                    when "0110100100" => data <= X"74";
                    when "0110100101" => data <= X"6f";
                    when "0110100110" => data <= X"20";
                    when "0110100111" => data <= X"00";
                    when "0110101000" => data <= X"0d";
                    when "0110101001" => data <= X"0a";
                    when "0110101010" => data <= X"45";
                    when "0110101011" => data <= X"52";
                    when "0110101100" => data <= X"52";
                    when "0110101101" => data <= X"4f";
                    when "0110101110" => data <= X"52";
                    when "0110101111" => data <= X"0d";
                    when "0110110000" => data <= X"0a";
                    when "0110110001" => data <= X"00";
                    when "0110110010" => data <= X"11";
                    when "0110110011" => data <= X"00";
                    when "0110110100" => data <= X"40";
                    when "0110110101" => data <= X"21";
                    when "0110110110" => data <= X"bf";
                    when "0110110111" => data <= X"01";
                    when "0110111000" => data <= X"01";
                    when "0110111001" => data <= X"4d";
                    when "0110111010" => data <= X"00";
                    when "0110111011" => data <= X"d5";
                    when "0110111100" => data <= X"ed";
                    when "0110111101" => data <= X"b0";
                    when "0110111110" => data <= X"c9";
                    when "0110111111" => data <= X"01";
                    when "0111000000" => data <= X"0c";
                    when "0111000001" => data <= X"bc";
                    when "0111000010" => data <= X"ed";
                    when "0111000011" => data <= X"49";
                    when "0111000100" => data <= X"01";
                    when "0111000101" => data <= X"30";
                    when "0111000110" => data <= X"bd";
                    when "0111000111" => data <= X"ed";
                    when "0111001000" => data <= X"49";
                    when "0111001001" => data <= X"21";
                    when "0111001010" => data <= X"00";
                    when "0111001011" => data <= X"c0";
                    when "0111001100" => data <= X"06";
                    when "0111001101" => data <= X"5a";
                    when "0111001110" => data <= X"af";
                    when "0111001111" => data <= X"70";
                    when "0111010000" => data <= X"23";
                    when "0111010001" => data <= X"bc";
                    when "0111010010" => data <= X"20";
                    when "0111010011" => data <= X"fb";
                    when "0111010100" => data <= X"01";
                    when "0111010101" => data <= X"81";
                    when "0111010110" => data <= X"7f";
                    when "0111010111" => data <= X"ed";
                    when "0111011000" => data <= X"49";
                    when "0111011001" => data <= X"01";
                    when "0111011010" => data <= X"fe";
                    when "0111011011" => data <= X"fe";
                    when "0111011100" => data <= X"3e";
                    when "0111011101" => data <= X"c0";
                    when "0111011110" => data <= X"ed";
                    when "0111011111" => data <= X"79";
                    when "0111100000" => data <= X"11";
                    when "0111100001" => data <= X"07";
                    when "0111100010" => data <= X"03";
                    when "0111100011" => data <= X"21";
                    when "0111100100" => data <= X"00";
                    when "0111100101" => data <= X"40";
                    when "0111100110" => data <= X"01";
                    when "0111100111" => data <= X"ff";
                    when "0111101000" => data <= X"fe";
                    when "0111101001" => data <= X"ed";
                    when "0111101010" => data <= X"49";
                    when "0111101011" => data <= X"ed";
                    when "0111101100" => data <= X"41";
                    when "0111101101" => data <= X"04";
                    when "0111101110" => data <= X"ed";
                    when "0111101111" => data <= X"51";
                    when "0111110000" => data <= X"ed";
                    when "0111110001" => data <= X"59";
                    when "0111110010" => data <= X"ed";
                    when "0111110011" => data <= X"61";
                    when "0111110100" => data <= X"ed";
                    when "0111110101" => data <= X"69";
                    when "0111110110" => data <= X"ed";
                    when "0111110111" => data <= X"78";
                    when "0111111000" => data <= X"3e";
                    when "0111111001" => data <= X"40";
                    when "0111111010" => data <= X"26";
                    when "0111111011" => data <= X"c0";
                    when "0111111100" => data <= X"ed";
                    when "0111111101" => data <= X"a2";
                    when "0111111110" => data <= X"04";
                    when "0111111111" => data <= X"bc";
                    when "1000000000" => data <= X"20";
                    when "1000000001" => data <= X"fa";
                    when "1000000010" => data <= X"05";
                    when "1000000011" => data <= X"ed";
                    when "1000000100" => data <= X"49";
                    when "1000000101" => data <= X"01";
                    when "1000000110" => data <= X"fe";
                    when "1000000111" => data <= X"fe";
                    when "1000001000" => data <= X"af";
                    when "1000001001" => data <= X"ed";
                    when "1000001010" => data <= X"79";
                    when "1000001011" => data <= X"c7";

	            when others => data <= X"00";
        	  end case;


    end process;

end impl;
